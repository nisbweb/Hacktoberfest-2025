// Design a 4-bit Carry Lookahead Adder using Verilog.

// The module should take two 4-bit inputs (A and B) and a carry-in.

// The outputs should be a 4-bit Sum and a carry-out.

// WRITE YOUR CODE HERE
