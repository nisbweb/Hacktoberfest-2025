// Design an Even Parity Generator for an 8-bit input using Verilog.

// The module should output a parity bit such that the total number of 1s

// (data + parity) is even.

// WRITE YOUR CODE HERE
