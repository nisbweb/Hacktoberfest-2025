// Design a BCD to 7-segment display decoder using Verilog.

// The module should take a 4-bit BCD input and generate outputs

// to drive a common cathode 7-segment display.

// WRITE YOUR CODE HERE
