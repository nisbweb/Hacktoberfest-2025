// Design a 4-bit Serial-In Parallel-Out (SIPO) Shift Register using Verilog.

// The module should take a serial input and shift data on every clock cycle.

// After 4 cycles, the output should be available in parallel (Q[3:0]).

// WRITE YOUR CODE HERE
